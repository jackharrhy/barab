module hello_world;

initial begin
  $display ("get barab'd");
  #10 $finish;
end

endmodule